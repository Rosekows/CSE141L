module lut_instr(
  input       [8:0] iptr,
  output logic[19:0] inst);
  always_comb begin case(iptr) 
    // product
    9'b000_000_000: inst = 20'b01110_00000_00000_00000; // done
    9'b000_000_001: inst = 20'b01100_00010_10001_00000; // ld	r2, [1]
    9'b000_000_010: inst = 20'b01100_00011_10010_00000; // ld 	r3, [2]	
    9'b000_000_011: inst = 20'b00011_00110_10001_00011; // and 	r6, 1, r3
    9'b000_000_100: inst = 20'b00110_00000_00000_00110; // cmp	r6, r0		// PSA: I changed the format of the compare instr
    9'b000_000_101: inst = 20'b00111_00000_00000_00100; // be	shift		// so they are now like:
    9'b000_000_110: inst = 20'b00000_00101_00010_00101; // add	r5, r2, r5	// [opcode] [00000] [in_b, either reg/constant] [in_a, reg]
    9'b000_000_111: inst = 20'b00000_00100_01000_00100; // add	r4, rO, r4  // Ex: cmp r7, r5 translates to opcode 00000 reg5 reg7
    9'b000_001_000: inst = 20'b00000_00100_00001_00100; // add 	r4, r1, r4	// and cmp r7, 10 translates to opcode 00000 constant10 reg7
    9'b000_001_001: inst = 20'b00011_00110_10011_00010; // and	r6, 128, r2
    9'b000_001_010: inst = 20'b00100_00010_10001_00010; // sll	r2, 1, r2
    9'b000_001_011: inst = 20'b00100_00001_10001_00001; // sll 	r1, 1, r1
    9'b000_001_100: inst = 20'b00000_00001_00110_00001; // add	r1, r6, r1
    9'b000_001_101: inst = 20'b00101_00011_10001_00011; // srl 	r3, 1, r3
    9'b000_001_110: inst = 20'b00000_00111_10001_00111; // add 	r7, 1, r7
    9'b000_001_111: inst = 20'b00110_00000_10100_00111; // cmp 	r7, 8
    9'b000_010_000: inst = 20'b01000_11111_11111_10011; // bl 	loop
    9'b000_010_001: inst = 20'b01001_00000_00000_00110; // bg 	lowerloop
    9'b000_010_010: inst = 20'b01100_00011_10101_00000; // ld	r3, [3]	
    9'b000_010_011: inst = 20'b01011_00010_00101_00000; // mov	r2, r5
    9'b000_010_100: inst = 20'b01011_00001_00100_00000; // mov 	r1, r4   
    
    9'b000_111_100: inst = 20'b01011_00101_00000_00000; // mov r5, r0
    9'b000_111_101: inst = 20'b01011_00100_00000_00000; // mov r4, r0
     
    9'b000_010_101: inst = 20'b00110_00000_11010_00111; // cmp	r7, 16   // so we don't have a 16 constant (can just add 1 and 15)
    9'b000_010_110: inst = 20'b01000_11111_11111_01011; // bl 	loop
    9'b000_010_111: inst = 20'b01101_00101_10111_00000; // st	[5], r5  // should this be st r5, [5]
    9'b000_011_000: inst = 20'b01101_00100_10110_00000; // st 	r4, [4]	

    // string match
    9'b000_011_001: inst = 20'b01100_00001_11000_00011; // ld	r1, [32 + r3]
    9'b000_011_010: inst = 20'b01100_00010_11001_00000; // ld 	r2, 6
    9'b000_011_011: inst = 20'b01011_00111_11010_00000; // mov	r7, 15
    9'b000_011_100: inst = 20'b00011_00110_00111_00001; // and	r6, r7, r1
    9'b000_011_101: inst = 20'b00010_00110_00010_00110; // xor	r6, r2, r6
    9'b000_011_110: inst = 20'b00110_00000_00000_00110; // cmp	r6, r0
    9'b000_011_111: inst = 20'b00111_00000_00000_00110; // be 	found
    9'b000_100_000: inst = 20'b00100_00111_10001_00111; // sll	r7, 1, r7
    9'b000_100_001: inst = 20'b00000_00100_10001_00100; // add 	r4, 1, r4
    9'b000_100_010: inst = 20'b00110_00000_10111_00100; // cmp 	r4, 5
    9'b000_100_011: inst = 20'b01000_11111_11111_11001; // bl	matchLoop
    9'b000_100_100: inst = 20'b01010_00000_00000_00010; // ba 	incJ
    9'b000_100_101: inst = 20'b00000_00101_10001_00101; // add	r5, 1, r5
    9'b000_100_110: inst = 20'b00000_00011_10001_00011; // add 	r3, 1, r3
    9'b000_100_111: inst = 20'b00110_00000_11011_00011; // cmp	r3, 64	
    9'b000_101_000: inst = 20'b01000_11111_11111_10001; // bl	stringLoop
    9'b000_101_001: inst = 20'b01101_00101_11100_00000; // st	r5, [7]

    // closest pair
    9'b000_101_010: inst = 20'b01011_00001_11101_00000; // mov	r1, 255
    9'b000_101_011: inst = 20'b01100_00100_10011_00010; // ld	r4, [128 + r2]
    9'b000_101_100: inst = 20'b00000_00011_10001_00010; // add	r3, 1, r2
    9'b000_101_101: inst = 20'b01100_00101_10011_00011; // ld	r5, [128 + r3]
    9'b000_101_110: inst = 20'b00110_00000_00101_00100; // cmp	r4, r5
    9'b000_101_111: inst = 20'b01001_00000_00000_00011; // bg	ijSub
    9'b000_110_000: inst = 20'b00001_00101_00101_00100; // sub	r5, r5, r4
    9'b000_110_001: inst = 20'b01010_00000_00000_00010; // ba	compDist
    9'b000_110_010: inst = 20'b00001_00101_00100_00101; // sub	r5, r4, r5
    9'b000_110_011: inst = 20'b00110_00000_00101_00001; // cmp	r1, r5
    9'b000_110_100: inst = 20'b01000_00000_00000_00010; // bl	incJ
    9'b000_110_101: inst = 20'b01011_00001_00101_00000; // mov	r1, r5
							// inc j
    9'b000_110_110: inst = 20'b00110_00000_11111_00011; // cmp	r3, 20
    9'b000_110_111: inst = 20'b01000_11111_11111_10101; // bl	inner
    9'b000_111_000: inst = 20'b00000_00010_10001_00010; // add 	r2, 1, r2
    9'b000_111_001: inst = 20'b00110_00000_11110_00010; // cmp	r2, 19
    9'b000_111_010: inst = 20'b01000_11111_11111_10000; // bl	outer
    9'b000_111_011: inst = 20'b01101_00001_10000_00000; // st	r1, [127]

    
    // MISC
    //9'b000_011_100: inst = 20'b01011_00111_11010_00000; // mov	r7, 15
    //9'b000_011_101: inst = 20'b01011_00001_11010_00000; // mov	r1, 15
    //9'b000_111_100: inst = 20'b00000_00111_10111_00111;  // add 	r7, 128, r7
    
  endcase
  //$display("Opcode is %d", inst[19:15]);
  end
endmodule